`include "mesi_coherency.v"

module mesi_coherency_tb ();

mesi_coherency dut (
);

endmodule
