// 8-way set associative cache
// cache replacement policy chosen is
// a 'least recently used' scheme
module l1cache_8w_sa (
);

endmodule
