// FSM based MESI protocol controller
module coherency_controller (
);

endmodule
