`include "l1cache_8w_sa.v"
`include "coherency_controller.v"

// top level block that comprises 4 L1 cache and
// snooping based MESI coherency controller
module mesi_coherency (
);

endmodule
